/*-----------------------------------------------------------------------------------------
MODULE FUNCTION :   Check the input signal (signal_in). Detects the presence of rising edge changes and output the result.
MODULE INPUT    : 
                    clk - clock signal of the current clock domain;
                    rst_n - reset signal of the module;
                    en - this makes the module work immediately
                    signal_in  - The signal (signal_in) be checked;
MODULE OUTPUT   :   
                    signal_out -   Outputs different values depending on the input signal;                          

AUTHOR               :   ljCai
MODIFICATION HISTORY :
VERSION     DATA            By           Change Description
---------------------------------------------------------------------------------------------
V0.1        23/01/16        ljCai       Original
V0.1        23/01/18        ljCai       Add enable signal; Synchronous Reset
-------------------------------------------------------------------------------------------*/
module rose (
    input   logic   clk         ,       //clock
    input   logic   rst_n       ,       //reset
    input   logic   en          ,       //enable signal
    input   logic   signal_in   ,       //input signal
    output  logic   match       ,       //match signal
    output  logic   fail                //fail signal
);
/*-------------------------------------------------------------
FUNCTION:Get the result of rose
-------------------------------------------------------------*/    
logic   delay_in_1  ;
logic   delay_in_2  ;
logic   en_1        ;
logic   en_2        ;   
always_ff @( posedge clk ) begin : rose_SV
        delay_in_1 <= signal_in ;
        delay_in_2 <= delay_in_1;
        en_1 <= en;
        en_2 <= en_1;
    if (rst_n == 1'b0) begin                //reset operation
        delay_in_1 <= 1'b0  ;
        delay_in_2 <= 1'b0  ;
    end
end
assign match = (~delay_in_2 & delay_in_1) & en_2 ;
assign fail  = ~match;
endmodule
//warning
